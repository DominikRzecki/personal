------------------------------------------------------------------------------------
--Project : DIC 4AHEL 
--Author  : Gr�bner
--Date    : 15/09/2020
--File    : DE10_Lite.vhd
--Design  : Terasic DE10 Board
------------------------------------------------------------------------------------
-- Description: Button Up/Down Counter, HEX
------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;

use work.DE10_Lite_const_pkg.ALL;

--=======================================================================================================
entity DE10_Lite is
  port (
        MAX10_CLK1_50 :  in std_logic;
        ---------------------------------------------------------------
        KEY           :  in std_logic_vector(    keys_c - 1 downto 0);
        SW            :  in std_logic_vector(switches_c - 1 downto 0);
        LEDR          : out std_logic_vector(    leds_c - 1 downto 0);
        ---------------------------------------------------------------
        HEX0          : out std_logic_vector(7 downto 0);
        HEX1          : out std_logic_vector(7 downto 0);
        HEX2          : out std_logic_vector(7 downto 0);
        HEX3          : out std_logic_vector(7 downto 0);
        HEX4          : out std_logic_vector(7 downto 0);
        HEX5          : out std_logic_vector(7 downto 0)
        ---------------------------------------------------------------
       );
end DE10_Lite;
--=======================================================================================================

--MAX10_CLK1_50 = not MAX10_CLK1_50 after de10_cycle_time_c;

architecture rtl of DE10_Lite is
  --=====================================================================================================
  
  --=====================================================================================================
begin
  --=====================================================================================================
  HEX0(7) <= '1';
  HEX1(7) <= '1';
  HEX2(7) <= '1';
  HEX3(7) <= '1';
  HEX4(7) <= '1';
  HEX5(7) <= '1';

  LEDR(1) <= not KEY(0);
  
  --=====================================================================================================
  BTN_1: entity work.debouncer(rtl)
  generic map (
    F_CLK => natural(de10_clk_freq_c),
    REQ_PRESS_TIME => 20 ms,
    SAMPLE_PERIOD => 500 us
  )
  port map (
    CLK => MAX10_CLK1_50,
    sig_in => KEY(0),
    sig_out => LEDR(0)
  );
  --=====================================================================================================

  --=====================================================================================================
end rtl;
--@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
